module top();


endmodule
