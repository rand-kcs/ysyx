module top(input a, input b, output f);

switch my_switch(a, b, f);

endmodule


