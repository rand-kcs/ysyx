module top(input clk, input rst, output [15:0] led);

light my_light(clk, rst, led);

endmodule
