module CSRs #(ADDR_WIDTH = 1, DATA_WIDTH = 1) (
  input clk,
  input rst,
  input valid_wbu,
  input [ADDR_WIDTH-1:0] waddr,
  input [DATA_WIDTH-1:0] wdata,
  //wen only stands for csrxx inst;
  input wen,
  input is_ecall_wbu,
  input is_mret_wbu,
  input [DATA_WIDTH-1:0] pc,

  input is_ecall_idu,
  input is_mret_idu,
  input [ADDR_WIDTH-1:0] raddr,
  output [DATA_WIDTH-1:0] data
);
// word_t mcause, mstatus, mepc;
// word_t mtvec;
/*
    case 0x300:
      return &(cpu.mstatus);
    case 0x305:
      return &(cpu.mtvec);
    case 0x341:
      return &(cpu.mepc);
    case 0x342:
      return &(cpu.mcause);
    case 0xF11:
      return &(cpu.mvendorid);
    case 0xF12:
      return &(cpu.marchid);
*/

reg [DATA_WIDTH-1:0] mcause;
reg [DATA_WIDTH-1:0] mstatus;

reg [DATA_WIDTH-1:0] mepc;
reg [DATA_WIDTH-1:0] mtvec;

reg [DATA_WIDTH-1:0] mvendorid;
reg [DATA_WIDTH-1:0] marchid;

wire [DATA_WIDTH-1:0] csr_data;

// WBU  control;
always@(posedge clk) begin
  if (rst) begin 
    mstatus <= 32'h1800;
    mvendorid <= 32'h79737978;
    marchid <= 32'd24100030;
  end
  if(valid_wbu) begin
    if(is_ecall_wbu) begin
      mepc <= pc;
      mcause  <= 32'hb;
    end
    else if(wen) begin
      case(waddr)
        12'h300: mstatus <= wdata; 
        12'h305: mtvec <= wdata; 
        12'h341: mepc <= wdata; 
        12'h342: mcause <= wdata;
        default: ;
      endcase
    end
  end
end


// IDU control
MuxKeyWithDefault #(6, 12, 32) csr_data_Mux(csr_data, raddr, 32'b0, {
  {12'h300} , mstatus,
  {12'h305} , mtvec ,
  {12'h341} , mepc ,
  {12'h342} , mcause,
  {12'hF11} , mvendorid ,
  {12'hF12} , marchid
});

wire [2:0] select;
assign select = {1'b0, is_ecall_idu, is_mret_idu};

MuxKeyWithDefault #(2, 3, 32) data_Mux(data, select, csr_data, {
  {3'b010}, mtvec,
  {3'b001}, mepc
});


endmodule
